------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 2.5
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : gtwizard_v2_5_gbe_gtx_exdes.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module gtwizard_v2_5_gbe_gtx_exdes
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_misc.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration************************

entity gtwizard_v2_5_gbe_gtx_exdes is
generic
(
    EXAMPLE_CONFIG_INDEPENDENT_LANES        : integer   := 1;
    EXAMPLE_LANE_WITH_START_CHAR            : integer   := 0;    -- specifies lane with unique start frame ch
    EXAMPLE_WORDS_IN_BRAM                   : integer   := 512;  -- specifies amount of data in BRAM
    EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "TRUE";    -- simulation setting for GT SecureIP model
    EXAMPLE_SIMULATION                      : integer   := 0;             -- Set to 1 for simulation
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 0           -- Set to 1 to use Chipscope to drive resets
);
port
(
    Q0_CLK1_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q0_CLK1_GTREFCLK_PAD_P_IN               : in   std_logic;
    DRP_CLK_IN                              : in   std_logic;
    SYSCLK_IN                               : in   std_logic;
    TRACK_DATA_OUT                          : out  std_logic;
    RXN_IN                                  : in   std_logic;
    RXP_IN                                  : in   std_logic;
    TXN_OUT                                 : out  std_logic;
    TXP_OUT                                 : out  std_logic
    
);


end gtwizard_v2_5_gbe_gtx_exdes;
    
architecture RTL of gtwizard_v2_5_gbe_gtx_exdes is

    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "gtwizard_v2_5_gbe_gtx,gtwizard_v2_5,{protocol_file=gigabit_ethernet_CC}";

--**************************Component Declarations*****************************


component gtwizard_v2_5_gbe_gtx_init 
generic
(
    -- Simulation attributes
    EXAMPLE_SIM_GTRESET_SPEEDUP    : string    := "FALSE";    -- Set to 1 to speed up sim reset
    EXAMPLE_SIMULATION             : integer   := 0;          -- Set to 1 for simulation
    EXAMPLE_USE_CHIPSCOPE          : integer   := 0           -- Set to 1 to use Chipscope to drive resets

);
port
(
    SYSCLK_IN                               : in   std_logic;
    SOFT_RESET_IN                           : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;

    --_________________________________________________________________________
    --GT0  (X1Y1)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT0_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT0_CPLLLOCK_OUT                        : out  std_logic;
    GT0_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT0_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT0_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT0_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT0_DRPCLK_IN                           : in   std_logic;
    GT0_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT0_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT0_DRPEN_IN                            : in   std_logic;
    GT0_DRPRDY_OUT                          : out  std_logic;
    GT0_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT0_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    GT0_RXPD_IN                             : in   std_logic_vector(1 downto 0);
    GT0_TXPD_IN                             : in   std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT0_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT0_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT0_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    GT0_RXCLKCORCNT_OUT                     : out  std_logic_vector(1 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT0_RXUSRCLK_IN                         : in   std_logic;
    GT0_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT0_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT0_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT0_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    GT0_GTXRXP_IN                           : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT0_GTXRXN_IN                           : in   std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    GT0_RXBUFRESET_IN                       : in   std_logic;
    GT0_RXBUFSTATUS_OUT                     : out  std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT0_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT0_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT0_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT0_GTRXRESET_IN                        : in   std_logic;
    GT0_RXPMARESET_IN                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    GT0_RXPOLARITY_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT0_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT0_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT0_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT0_GTTXRESET_IN                        : in   std_logic;
    GT0_TXUSERRDY_IN                        : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    GT0_TXCHARDISPMODE_IN                   : in   std_logic_vector(1 downto 0);
    GT0_TXCHARDISPVAL_IN                    : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT0_TXUSRCLK_IN                         : in   std_logic;
    GT0_TXUSRCLK2_IN                        : in   std_logic;
    --------------------- Transmit Ports - PCI Express Ports -------------------
    GT0_TXELECIDLE_IN                       : in   std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    GT0_TXBUFSTATUS_OUT                     : out  std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT0_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT0_GTXTXN_OUT                          : out  std_logic;
    GT0_GTXTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT0_TXOUTCLK_OUT                        : out  std_logic;
    GT0_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT0_TXOUTCLKPCS_OUT                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    GT0_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT0_TXRESETDONE_OUT                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    GT0_TXPOLARITY_IN                       : in   std_logic;
   

    --____________________________COMMON PORTS________________________________
    ---------------------- Common Block  - Ref Clock Ports ---------------------
    GT0_GTREFCLK0_COMMON_IN                 : in   std_logic;
    ------------------------- Common Block - QPLL Ports ------------------------
    GT0_QPLLLOCK_OUT                        : out  std_logic;
    GT0_QPLLLOCKDETCLK_IN                   : in   std_logic;
    GT0_QPLLRESET_IN                        : in   std_logic


);
end component;

component gtwizard_v2_5_gbe_gtx_GT_USRCLK_SOURCE 
port
(
    Q0_CLK1_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q0_CLK1_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q0_CLK1_GTREFCLK_OUT                    : out  std_logic;
 
    GT0_TXUSRCLK_OUT             : out std_logic;
    GT0_TXUSRCLK2_OUT            : out std_logic;
    GT0_TXOUTCLK_IN              : in  std_logic;
    GT0_RXUSRCLK_OUT             : out std_logic;
    GT0_RXUSRCLK2_OUT            : out std_logic;
    GT0_RXOUTCLK_IN              : in  std_logic;
    DRPCLK_IN                          : in  std_logic;
    DRPCLK_OUT                         : out std_logic
);
end component;




component gtwizard_v2_5_gbe_gtx_GT_FRAME_GEN 
generic
(
     WORDS_IN_BRAM    : integer := 512
);
port
(
    -- User Interface
    TX_DATA_OUT             : out   std_logic_vector(79 downto 0);
    TXCTRL_OUT              : out   std_logic_vector(7 downto 0); 
    -- System Interface
    USER_CLK                : in    std_logic;      
    SYSTEM_RESET            : in    std_logic
); 
end component;

component gtwizard_v2_5_gbe_gtx_GT_FRAME_CHECK 
generic
(
    RX_DATA_WIDTH            : integer := 16;
    RXCTRL_WIDTH             : integer := 2; 
    WORDS_IN_BRAM            : integer := 256;
    CHANBOND_SEQ_LEN         : integer := 1;
    COMMA_DOUBLE             : std_logic_vector(15 downto 0) := x"f628";
    START_OF_PACKET_CHAR     : std_logic_vector(15 downto 0) := x"02bc"
);
port
(
    -- User Interface
    RX_DATA_IN               : in  std_logic_vector((RX_DATA_WIDTH-1) downto 0);
    RXCTRL_IN                : in  std_logic_vector((RXCTRL_WIDTH-1) downto 0); 
    RXENMCOMMADET_OUT        : out std_logic;
    RXENPCOMMADET_OUT        : out std_logic;
    RX_ENCHAN_SYNC_OUT       : out std_logic;
    RX_CHANBOND_SEQ_IN       : in  std_logic;

    -- Control Interface
    INC_IN                   : in  std_logic; 
    INC_OUT                  : out std_logic; 
    PATTERN_MATCHB_OUT       : out std_logic;
    RESET_ON_ERROR_IN        : in  std_logic;


    -- Error Monitoring
    ERROR_COUNT_OUT          : out std_logic_vector(7 downto 0);

    -- Track Data
    TRACK_DATA_OUT           : out std_logic;

 

    -- System Interface
    USER_CLK                 : in std_logic;       
    SYSTEM_RESET             : in std_logic
);
end component;

-- Chipscope modules
attribute syn_black_box                : boolean;
attribute syn_noprune                  : boolean;


component data_vio
port
(
    control                 : inout std_logic_vector(35 downto 0);
    clk                     : in    std_logic;
    async_in                : in    std_logic_vector(31 downto 0);
    async_out               : out   std_logic_vector(31 downto 0);
    sync_in                 : in    std_logic_vector(31 downto 0);
    sync_out                : out   std_logic_vector(31 downto 0)
);
end component;
attribute syn_black_box of data_vio : component is TRUE;
attribute syn_noprune of data_vio   : component is TRUE;


component icon
port
(
    control0                : inout std_logic_vector(35 downto 0);
    control1                : inout std_logic_vector(35 downto 0);
    control2                : inout std_logic_vector(35 downto 0);
    control3                : inout std_logic_vector(35 downto 0);
    control4                : inout std_logic_vector(35 downto 0);
    control5                : inout std_logic_vector(35 downto 0)
);
end component;
attribute syn_black_box of icon : component is TRUE;
attribute syn_noprune of icon   : component is TRUE;


component ila
port
(
    control                 : inout std_logic_vector(35 downto 0);
    clk                     : in    std_logic;
    trig0                   : in    std_logic_vector(163 downto 0)
);
end component;

--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--************************** Register Declarations ****************************

    signal   gt0_txfsmresetdone_i            : std_logic;
    signal   gt0_rxfsmresetdone_i            : std_logic;
    signal   gt0_txfsmresetdone_r            : std_logic;
    signal   gt0_txfsmresetdone_r2           : std_logic;
    signal   gt0_rxresetdone_r               : std_logic;
    signal   gt0_rxresetdone_r2              : std_logic;
    signal   gt0_rxresetdone_r3              : std_logic;


    signal   reset_pulse                     : std_logic_vector(3 downto 0);
    signal   reset_counter  :   unsigned(5 downto 0) := "000000";


--**************************** Wire Declarations ******************************
    -------------------------- GT Wrapper Wires ------------------------------
    --________________________________________________________________________
    --________________________________________________________________________
    --GT0   (X1Y1)

    --------------------------------- CPLL Ports -------------------------------
    signal  gt0_cpllfbclklost_i             : std_logic;
    signal  gt0_cplllock_i                  : std_logic;
    signal  gt0_cpllrefclklost_i            : std_logic;
    signal  gt0_cpllreset_i                 : std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt0_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt0_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt0_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt0_drpen_i                     : std_logic;
    signal  gt0_drprdy_i                    : std_logic;
    signal  gt0_drpwe_i                     : std_logic;
    ------------------------------- Loopback Ports -----------------------------
    signal  gt0_loopback_i                  : std_logic_vector(2 downto 0);
    ------------------------------ Power-Down Ports ----------------------------
    signal  gt0_rxpd_i                      : std_logic_vector(1 downto 0);
    signal  gt0_txpd_i                      : std_logic_vector(1 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt0_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt0_eyescandataerror_i          : std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    signal  gt0_rxcdrlock_i                 : std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    signal  gt0_rxclkcorcnt_i               : std_logic_vector(1 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt0_rxdata_i                    : std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt0_rxdisperr_i                 : std_logic_vector(1 downto 0);
    signal  gt0_rxnotintable_i              : std_logic_vector(1 downto 0);
    --------------------------- Receive Ports - RX AFE -------------------------
    signal  gt0_gtxrxp_i                    : std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt0_gtxrxn_i                    : std_logic;
    ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
    signal  gt0_rxbufreset_i                : std_logic;
    signal  gt0_rxbufstatus_i               : std_logic_vector(2 downto 0);
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt0_rxmcommaalignen_i           : std_logic;
    signal  gt0_rxpcommaalignen_i           : std_logic;
    --------------------- Receive Ports - RX Equilizer Ports -------------------
    signal  gt0_rxlpmhfhold_i               : std_logic;
    signal  gt0_rxlpmlfhold_i               : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt0_rxoutclk_i                  : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt0_gtrxreset_i                 : std_logic;
    signal  gt0_rxpcsreset_i                : std_logic;
    signal  gt0_rxpmareset_i                : std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    signal  gt0_rxpolarity_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt0_rxchariscomma_i             : std_logic_vector(1 downto 0);
    signal  gt0_rxcharisk_i                 : std_logic_vector(1 downto 0);
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt0_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt0_gttxreset_i                 : std_logic;
    signal  gt0_txuserrdy_i                 : std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    signal  gt0_txchardispmode_i            : std_logic_vector(1 downto 0);
    signal  gt0_txchardispval_i             : std_logic_vector(1 downto 0);
    --------------------- Transmit Ports - PCI Express Ports -------------------
    signal  gt0_txelecidle_i                : std_logic;
    ---------------------- Transmit Ports - TX Buffer Ports --------------------
    signal  gt0_txbufstatus_i               : std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt0_txdata_i                    : std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt0_gtxtxn_i                    : std_logic;
    signal  gt0_gtxtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt0_txoutclk_i                  : std_logic;
    signal  gt0_txoutclkfabric_i            : std_logic;
    signal  gt0_txoutclkpcs_i               : std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    signal  gt0_txcharisk_i                 : std_logic_vector(1 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt0_txpcsreset_i                : std_logic;
    signal  gt0_txresetdone_i               : std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    signal  gt0_txpolarity_i                : std_logic;



    --____________________________COMMON PORTS________________________________
    ------------------------- Common Block - QPLL Ports ------------------------
    signal  gt0_qplllock_i                  : std_logic;
    signal  gt0_qpllrefclklost_i            : std_logic;
    signal  gt0_qpllreset_i                 : std_logic;



    ------------------------------- Global Signals -----------------------------
    signal  gt0_tx_system_reset_c           : std_logic;
    signal  gt0_rx_system_reset_c           : std_logic;
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_ground_vec_i            : std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   : std_logic;
    signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
    signal  drpclk_in_i                     : std_logic;
 
    signal  GTTXRESET_IN                    : std_logic;
    signal  GTRXRESET_IN                    : std_logic;
    signal  CPLLRESET_IN                    : std_logic;
    signal  QPLLRESET_IN                    : std_logic;

   ------------------------------- User Clocks ---------------------------------
    attribute keep: string;
    signal    gt0_txusrclk_i                  : std_logic; 
    signal    gt0_txusrclk2_i                 : std_logic; 
    signal    gt0_rxusrclk_i                  : std_logic; 
    signal    gt0_rxusrclk2_i                 : std_logic; 
    attribute keep of gt0_txusrclk_i : signal is "true";
    attribute keep of gt0_txusrclk2_i : signal is "true";
    attribute keep of gt0_rxusrclk_i : signal is "true";
    attribute keep of gt0_rxusrclk2_i : signal is "true";
 

    ----------------------------- Reference Clocks ----------------------------
    
    signal    q0_clk1_refclk_i                : std_logic;


    ----------------------- Frame check/gen Module Signals --------------------
    
    signal    gt0_matchn_i                    : std_logic;
    
    signal    gt0_txcharisk_float_i           : std_logic_vector(5 downto 0);
    
    signal    gt0_txdata_float16_i            : std_logic_vector(15 downto 0);
    signal    gt0_txdata_float_i              : std_logic_vector(47 downto 0);
    
    signal    gt0_track_data_i                : std_logic;
    signal    gt0_block_sync_i                : std_logic;
    signal    gt0_error_count_i               : std_logic_vector(7 downto 0);
    signal    gt0_frame_check_reset_i         : std_logic;
    signal    gt0_inc_in_i                    : std_logic;
    signal    gt0_inc_out_i                   : std_logic;
    signal    gt0_unscrambled_data_i          : std_logic_vector(15 downto 0);

    signal    reset_on_data_error_i           : std_logic;
    signal    track_data_out_i                : std_logic;
   

    ----------------------- Chipscope Signals ---------------------------------

    signal  tx_data_vio_control_i           : std_logic_vector(35 downto 0);
    signal  rx_data_vio_control_i           : std_logic_vector(35 downto 0);
    signal  shared_vio_control_i            : std_logic_vector(35 downto 0);
    signal  ila_control_i                   : std_logic_vector(35 downto 0);
    signal  channel_drp_vio_control_i       : std_logic_vector(35 downto 0);
    signal  common_drp_vio_control_i        : std_logic_vector(35 downto 0);
    signal  tx_data_vio_async_in_i          : std_logic_vector(31 downto 0);
    signal  tx_data_vio_sync_in_i           : std_logic_vector(31 downto 0);
    signal  tx_data_vio_async_out_i         : std_logic_vector(31 downto 0);
    signal  tx_data_vio_sync_out_i          : std_logic_vector(31 downto 0);
    signal  rx_data_vio_async_in_i          : std_logic_vector(31 downto 0);
    signal  rx_data_vio_sync_in_i           : std_logic_vector(31 downto 0);
    signal  rx_data_vio_async_out_i         : std_logic_vector(31 downto 0);
    signal  rx_data_vio_sync_out_i          : std_logic_vector(31 downto 0);
    signal  shared_vio_in_i                 : std_logic_vector(31 downto 0);
    signal  shared_vio_out_i                : std_logic_vector(31 downto 0);
    signal  ila_in_i                        : std_logic_vector(163 downto 0);
    signal  channel_drp_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  channel_drp_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  channel_drp_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  channel_drp_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  common_drp_vio_async_in_i       : std_logic_vector(31 downto 0);
    signal  common_drp_vio_sync_in_i        : std_logic_vector(31 downto 0);
    signal  common_drp_vio_async_out_i      : std_logic_vector(31 downto 0);
    signal  common_drp_vio_sync_out_i       : std_logic_vector(31 downto 0);

    signal  gt0_tx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt0_tx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt0_tx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt0_tx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt0_rx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt0_rx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt0_rx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt0_rx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt0_ila_in_i                    : std_logic_vector(163 downto 0);
    signal  gt0_channel_drp_vio_async_in_i  : std_logic_vector(31 downto 0);
    signal  gt0_channel_drp_vio_sync_in_i   : std_logic_vector(31 downto 0);
    signal  gt0_channel_drp_vio_async_out_i : std_logic_vector(31 downto 0);
    signal  gt0_channel_drp_vio_sync_out_i  : std_logic_vector(31 downto 0);
    signal  gt0_common_drp_vio_async_in_i   : std_logic_vector(31 downto 0);
    signal  gt0_common_drp_vio_sync_in_i    : std_logic_vector(31 downto 0);
    signal  gt0_common_drp_vio_async_out_i  : std_logic_vector(31 downto 0);
    signal  gt0_common_drp_vio_sync_out_i   : std_logic_vector(31 downto 0);


    signal    gttxreset_i                     : std_logic;
    signal    gtrxreset_i                     : std_logic;

    signal    user_tx_reset_i                 : std_logic;
    signal    user_rx_reset_i                 : std_logic;
    signal    tx_vio_clk_i                    : std_logic;
    signal    tx_vio_clk_mux_out_i            : std_logic;    
    signal    rx_vio_ila_clk_i                : std_logic;
    signal    rx_vio_ila_clk_mux_out_i        : std_logic;    

    
    signal    cpllreset_i                     : std_logic;
    


   function and_reduce(arg: std_logic_vector) return std_logic is
	variable result: std_logic;
    begin
	result := '1';
	for i in arg'range loop
	    result := result and arg(i);
	end loop;
        return result;
    end;


--**************************** Main Body of Code *******************************
begin

    --  Static signal Assigments
    tied_to_ground_i                             <= '0';
    tied_to_ground_vec_i                         <= x"0000000000000000";
    tied_to_vcc_i                                <= '1';
    tied_to_vcc_vec_i                            <= x"ff";

    
  
    gt0_usrclk_source : gtwizard_v2_5_gbe_gtx_GT_USRCLK_SOURCE
    port map
    (
        Q0_CLK1_GTREFCLK_PAD_N_IN       =>      Q0_CLK1_GTREFCLK_PAD_N_IN,
        Q0_CLK1_GTREFCLK_PAD_P_IN       =>      Q0_CLK1_GTREFCLK_PAD_P_IN,
        Q0_CLK1_GTREFCLK_OUT            =>      q0_clk1_refclk_i,
 
        GT0_TXUSRCLK_OUT                =>      gt0_txusrclk_i,
        GT0_TXUSRCLK2_OUT               =>      gt0_txusrclk2_i,
        GT0_TXOUTCLK_IN                 =>      gt0_txoutclk_i,
        GT0_RXUSRCLK_OUT                =>      gt0_rxusrclk_i,
        GT0_RXUSRCLK2_OUT               =>      gt0_rxusrclk2_i,
        GT0_RXOUTCLK_IN                 =>      gt0_rxoutclk_i,
        DRPCLK_IN                       =>      DRP_CLK_IN,
        DRPCLK_OUT                      =>      drpclk_in_i

    );


    ----------------------------- The GT Wrapper -----------------------------
    
    -- Use the instantiation template in the example directory to add the GT wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.


    gtwizard_v2_5_gbe_gtx_init_i : gtwizard_v2_5_gbe_gtx_init
    generic map
    (
        EXAMPLE_SIM_GTRESET_SPEEDUP     =>      EXAMPLE_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION              =>      EXAMPLE_SIMULATION,
        EXAMPLE_USE_CHIPSCOPE           =>      EXAMPLE_USE_CHIPSCOPE
    )
    port map
    (
        SYSCLK_IN                       =>      SYSCLK_IN,
        SOFT_RESET_IN                   =>      tied_to_ground_i,
        DONT_RESET_ON_DATA_ERROR_IN     =>      tied_to_ground_i,
        GT0_TX_FSM_RESET_DONE_OUT       =>      gt0_txfsmresetdone_i,
        GT0_RX_FSM_RESET_DONE_OUT       =>      gt0_rxfsmresetdone_i,
        GT0_DATA_VALID_IN               =>      gt0_track_data_i,

  
 
 
 
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT0  (X1Y1)

        --------------------------------- CPLL Ports -------------------------------
        GT0_CPLLFBCLKLOST_OUT           =>      gt0_cpllfbclklost_i,
        GT0_CPLLLOCK_OUT                =>      gt0_cplllock_i,
        GT0_CPLLLOCKDETCLK_IN           =>      drpclk_in_i,
        GT0_CPLLRESET_IN                =>      gt0_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        GT0_GTREFCLK0_IN                =>      q0_clk1_refclk_i,
        ---------------------------- Channel - DRP Ports  --------------------------
        GT0_DRPADDR_IN                  =>      gt0_drpaddr_i,
        GT0_DRPCLK_IN                   =>      drpclk_in_i,
        GT0_DRPDI_IN                    =>      gt0_drpdi_i,
        GT0_DRPDO_OUT                   =>      gt0_drpdo_i,
        GT0_DRPEN_IN                    =>      gt0_drpen_i,
        GT0_DRPRDY_OUT                  =>      gt0_drprdy_i,
        GT0_DRPWE_IN                    =>      gt0_drpwe_i,
        ------------------------------- Loopback Ports -----------------------------
        GT0_LOOPBACK_IN                 =>      "000",
        ------------------------------ Power-Down Ports ----------------------------
        GT0_RXPD_IN                     =>      gt0_rxpd_i,
        GT0_TXPD_IN                     =>      gt0_txpd_i,
        --------------------- RX Initialization and Reset Ports --------------------
        GT0_RXUSERRDY_IN                =>      gt0_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        GT0_EYESCANDATAERROR_OUT        =>      gt0_eyescandataerror_i,
        ------------------------- Receive Ports - CDR Ports ------------------------
        GT0_RXCDRLOCK_OUT               =>      gt0_rxcdrlock_i,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        GT0_RXCLKCORCNT_OUT             =>      gt0_rxclkcorcnt_i,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        GT0_RXUSRCLK_IN                 =>      gt0_rxusrclk_i,
        GT0_RXUSRCLK2_IN                =>      gt0_rxusrclk_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        GT0_RXDATA_OUT                  =>      gt0_rxdata_i,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        GT0_RXDISPERR_OUT               =>      gt0_rxdisperr_i,
        GT0_RXNOTINTABLE_OUT            =>      gt0_rxnotintable_i,
        --------------------------- Receive Ports - RX AFE -------------------------
        GT0_GTXRXP_IN                   =>      RXP_IN,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GT0_GTXRXN_IN                   =>      RXN_IN,
        ------------------- Receive Ports - RX Buffer Bypass Ports -----------------
        GT0_RXBUFRESET_IN               =>      gt0_rxbufreset_i,
        GT0_RXBUFSTATUS_OUT             =>      gt0_rxbufstatus_i,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        GT0_RXMCOMMAALIGNEN_IN          =>      gt0_rxmcommaalignen_i,
        GT0_RXPCOMMAALIGNEN_IN          =>      gt0_rxpcommaalignen_i,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        GT0_RXOUTCLK_OUT                =>      gt0_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GT0_GTRXRESET_IN                =>      gt0_gtrxreset_i,
        GT0_RXPMARESET_IN               =>      gt0_rxpmareset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        GT0_RXPOLARITY_IN               =>      gt0_rxpolarity_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        GT0_RXCHARISCOMMA_OUT           =>      gt0_rxchariscomma_i,
        GT0_RXCHARISK_OUT               =>      gt0_rxcharisk_i,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        GT0_RXRESETDONE_OUT             =>      gt0_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        GT0_GTTXRESET_IN                =>      gt0_gttxreset_i,
        GT0_TXUSERRDY_IN                =>      gt0_txuserrdy_i,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        GT0_TXCHARDISPMODE_IN           =>      gt0_txchardispmode_i,
        GT0_TXCHARDISPVAL_IN            =>      gt0_txchardispval_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        GT0_TXUSRCLK_IN                 =>      gt0_txusrclk_i,
        GT0_TXUSRCLK2_IN                =>      gt0_txusrclk_i,
        --------------------- Transmit Ports - PCI Express Ports -------------------
        GT0_TXELECIDLE_IN               =>      gt0_txelecidle_i,
        ---------------------- Transmit Ports - TX Buffer Ports --------------------
        GT0_TXBUFSTATUS_OUT             =>      gt0_txbufstatus_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        GT0_TXDATA_IN                   =>      gt0_txdata_i,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GT0_GTXTXN_OUT                  =>      TXN_OUT,
        GT0_GTXTXP_OUT                  =>      TXP_OUT,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        GT0_TXOUTCLK_OUT                =>      gt0_txoutclk_i,
        GT0_TXOUTCLKFABRIC_OUT          =>      gt0_txoutclkfabric_i,
        GT0_TXOUTCLKPCS_OUT             =>      gt0_txoutclkpcs_i,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        GT0_TXCHARISK_IN                =>      gt0_txcharisk_i,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        GT0_TXRESETDONE_OUT             =>      gt0_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        GT0_TXPOLARITY_IN               =>      gt0_txpolarity_i,




    --____________________________COMMON PORTS________________________________
        ---------------------- Common Block  - Ref Clock Ports ---------------------
        GT0_GTREFCLK0_COMMON_IN         =>      q0_clk1_refclk_i,
        ------------------------- Common Block - QPLL Ports ------------------------
        GT0_QPLLLOCK_OUT                =>      gt0_qplllock_i,
        GT0_QPLLLOCKDETCLK_IN           =>      drpclk_in_i,
        GT0_QPLLRESET_IN                =>      gt0_qpllreset_i

    );



    -------------------------- User Module Resets -----------------------------
    -- All the User Modules i.e. FRAME_GEN, FRAME_CHECK and the sync modules
    -- are held in reset till the RESETDONE goes high. 
    -- The RESETDONE is registered a couple of times on USRCLK2 and connected 
    -- to the reset of the modules
    
    process( gt0_rxusrclk_i,gt0_rxresetdone_i)
    begin
        if(gt0_rxresetdone_i = '0') then
            gt0_rxresetdone_r  <= '0'   after DLY;
            gt0_rxresetdone_r2 <= '0'   after DLY;
            gt0_rxresetdone_r3 <= '0'   after DLY;
        elsif(gt0_rxusrclk_i'event and gt0_rxusrclk_i = '1') then
            gt0_rxresetdone_r  <= gt0_rxresetdone_i   after DLY;
            gt0_rxresetdone_r2 <= gt0_rxresetdone_r   after DLY;
            gt0_rxresetdone_r3  <= gt0_rxresetdone_r2   after DLY;
        end if;
    end process;

    process( gt0_txusrclk_i,gt0_txfsmresetdone_i)
    begin
        if(gt0_txfsmresetdone_i = '0') then
            gt0_txfsmresetdone_r  <= '0'   after DLY;
            gt0_txfsmresetdone_r2 <= '0'   after DLY;
        elsif(gt0_txusrclk_i'event and gt0_txusrclk_i = '1') then
            gt0_txfsmresetdone_r  <= gt0_txfsmresetdone_i   after DLY;
            gt0_txfsmresetdone_r2 <= gt0_txfsmresetdone_r   after DLY;
        end if;
    end process;

    ------------------------------ Frame Generators ---------------------------
    -- The example design uses Block RAM based frame generators to provide test
    -- data to the GTs for transmission. By default the frame generators are 
    -- loaded with an incrementing data sequence that includes commas/alignment
    -- characters for alignment. If your protocol uses channel bonding, the 
    -- frame generator will also be preloaded with a channel bonding sequence.
    
    -- You can modify the data transmitted by changing the INIT values of the frame
    -- generator in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.

    gt0_frame_gen : gtwizard_v2_5_gbe_gtx_GT_FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM
    )
    port map
    (
        -- User Interface
        TX_DATA_OUT(79 downto 32)       =>      gt0_txdata_float_i,
        TX_DATA_OUT(15 downto 0)        =>      gt0_txdata_float16_i,
        TX_DATA_OUT(31 downto 16)       =>      gt0_txdata_i,
 
        TXCTRL_OUT(7 downto 2)          =>      gt0_txcharisk_float_i,
        TXCTRL_OUT(1 downto 0)          =>      gt0_txcharisk_i,
        -- System Interface
        USER_CLK                        =>      gt0_txusrclk_i,
        SYSTEM_RESET                    =>      gt0_tx_system_reset_c
    );
    


    ---------------------------------- Frame Checkers -------------------------
    -- The example design uses Block RAM based frame checkers to verify incoming  
    -- data. By default the frame generators are loaded with a data sequence that 
    -- matches the outgoing sequence of the frame generators for the TX ports.
    
    -- You can modify the expected data sequence by changing the INIT values of the frame
    -- checkers in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.
    
    -- When the frame checker receives data, it attempts to synchronise to the 
    -- incoming pattern by looking for the first sequence in the pattern. Once it 
    -- finds the first sequence, it increments through the sequence, and indicates an 
    -- error whenever the next value received does not match the expected value.

    gt0_frame_check_reset_i                      <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else gt0_matchn_i;

    -- gt0_frame_check0 is always connected to the lane with the start of char
    -- and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
    gt0_inc_in_i                                 <= '0';

    gt0_frame_check : gtwizard_v2_5_gbe_gtx_GT_FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      16,
        RXCTRL_WIDTH                    =>      2,
        COMMA_DOUBLE                    =>      x"02bc",
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        START_OF_PACKET_CHAR            =>      x"02bc"
    )
    port map
    (
        -- GT Interface
        RX_DATA_IN                      =>      gt0_rxdata_i,
        RXCTRL_IN                       =>      gt0_rxcharisk_i,
        RXENMCOMMADET_OUT               =>      gt0_rxmcommaalignen_i,
        RXENPCOMMADET_OUT               =>      gt0_rxpcommaalignen_i,
        RX_ENCHAN_SYNC_OUT              =>      open,
        RX_CHANBOND_SEQ_IN              =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      gt0_inc_in_i,
        INC_OUT                         =>      gt0_inc_out_i,
        PATTERN_MATCHB_OUT              =>      gt0_matchn_i,
        RESET_ON_ERROR_IN               =>      gt0_frame_check_reset_i,
        -- System Interface
        USER_CLK                        =>      gt0_rxusrclk_i,
        SYSTEM_RESET                    =>      gt0_rx_system_reset_c,
        ERROR_COUNT_OUT                 =>      gt0_error_count_i,
        TRACK_DATA_OUT                  =>      gt0_track_data_i
    );




    TRACK_DATA_OUT                               <= track_data_out_i;

    track_data_out_i                             <= 
                                gt0_track_data_i ;








-------------------------------------------------------------------------------
    
    
    
    
    

----------------------------- Chipscope Connections -----------------------
    -- When the example design is run in hardware, it uses chipscope to allow the
    -- example design and GT wrapper to be controlled and monitored. The 
    -- EXAMPLE_USE_CHIPSCOPE parameter allows chipscope to be removed for simulation.

chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate
    
    -- ICON for all VIOs 
    icon_i : icon
    port map
    (
        control0                        =>      shared_vio_control_i,
        control1                        =>      tx_data_vio_control_i,
        control2                        =>      rx_data_vio_control_i,
        control3                        =>      ila_control_i,
        control4                        =>      channel_drp_vio_control_i,
        control5                        =>      common_drp_vio_control_i
    );

    -- Shared VIO for Channel DRP  
    channel_drp_i : data_vio 
    port map
    (
        control                         =>      channel_drp_vio_control_i,
        async_in                        =>      channel_drp_vio_async_in_i,
        async_out                       =>      channel_drp_vio_async_out_i,
        sync_in                         =>      channel_drp_vio_sync_in_i,
        sync_out                        =>      channel_drp_vio_sync_out_i,
        clk                             =>      drpclk_in_i
    );

    -- Shared VIO for Quad common DRP  
    common_drp_i : data_vio 
    port map
    (
        control                         =>      common_drp_vio_control_i,
        async_in                        =>      common_drp_vio_async_in_i,
        async_out                       =>      common_drp_vio_async_out_i,
        sync_in                         =>      common_drp_vio_sync_in_i,
        sync_out                        =>      common_drp_vio_sync_out_i,
        clk                             =>      drpclk_in_i
    );

    -- Shared VIO for all transievers 
    shared_vio_i : data_vio
    port map
    (
        control                         =>      shared_vio_control_i,
        clk                             =>      tied_to_ground_i,
        async_in                        =>      shared_vio_in_i,
        async_out                       =>      shared_vio_out_i,
        sync_in                         =>      tied_to_ground_vec_i(31 downto 0),
        sync_out                        =>      open
    );
    
    
    -- TX VIO 
    tx_data_vio_i : data_vio
    port map
    (
        control                         =>      tx_data_vio_control_i,
        clk                             =>      gt0_txusrclk_i,
        async_in                        =>      tx_data_vio_async_in_i,
        async_out                       =>      tx_data_vio_async_out_i,
        sync_in                         =>      tx_data_vio_sync_in_i,
        sync_out                        =>      tx_data_vio_sync_out_i
    );
    
    -- RX VIO 
    rx_data_vio_i : data_vio
    port map
    (
        control                         =>      rx_data_vio_control_i,
        clk                             =>      gt0_rxusrclk_i,
        async_in                        =>      rx_data_vio_async_in_i,
        async_out                       =>      rx_data_vio_async_out_i,
        sync_in                         =>      rx_data_vio_sync_in_i,
        sync_out                        =>      rx_data_vio_sync_out_i
    );
    
    -- RX ILA
    ila_i : ila
    port map
    (
        control                         =>      ila_control_i,
        clk                             =>      gt0_rxusrclk_i,
        trig0                           =>      ila_in_i
    );



    -- assign resets for frame_gen modules
    gt0_tx_system_reset_c                        <= not gt0_txfsmresetdone_r2 or user_tx_reset_i;

    -- assign resets for frame_check modules
    gt0_rx_system_reset_c                        <= not gt0_rxresetdone_r3 or user_rx_reset_i;

    gt0_gtrxreset_i                              <= gtrxreset_i or not gt0_cplllock_i;
    gt0_gttxreset_i                              <= gttxreset_i or not gt0_cplllock_i;

    gt0_cpllreset_i                              <= cpllreset_i;


    -- Shared VIO Outputs
    gttxreset_i                                  <= shared_vio_out_i(31);
    gtrxreset_i                                  <= shared_vio_out_i(30);
    user_tx_reset_i                              <= shared_vio_out_i(29);
    user_rx_reset_i                              <= shared_vio_out_i(28);
    cpllreset_i                                  <= shared_vio_out_i(27);

    -- Shared VIO Inputs
    shared_vio_in_i(31 downto 0)                 <= "00000000000000000000000000000000";

    -- Chipscope connections on GT 0
    gt0_tx_data_vio_async_in_i(31 downto 0)      <= "00000000000000000000000000000000";
    gt0_tx_data_vio_sync_in_i(31)                <= gt0_txresetdone_i;
    gt0_tx_data_vio_sync_in_i(30 downto 29)      <= gt0_txbufstatus_i;
    gt0_tx_data_vio_sync_in_i(28 downto 0)       <= "00000000000000000000000000000";
    gt0_loopback_i                               <= tx_data_vio_async_out_i(31 downto 29);
    gt0_txuserrdy_i                              <= tx_data_vio_sync_out_i(31);
    gt0_txpd_i                                   <= tx_data_vio_sync_out_i(30 downto 29);
    gt0_txchardispmode_i                         <= tx_data_vio_sync_out_i(28 downto 27);
    gt0_txchardispval_i                          <= tx_data_vio_sync_out_i(26 downto 25);
    gt0_txpolarity_i                             <= tx_data_vio_sync_out_i(24);
    gt0_txelecidle_i                             <= tx_data_vio_sync_out_i(23);
    gt0_rx_data_vio_async_in_i(31 downto 0)      <= "00000000000000000000000000000000";
    gt0_rx_data_vio_sync_in_i(31)                <= gt0_rxresetdone_i;
    gt0_rx_data_vio_sync_in_i(30 downto 0)       <= "0000000000000000000000000000000";
    gt0_rxuserrdy_i                              <= rx_data_vio_async_out_i(31);
    gt0_rxpd_i                                   <= rx_data_vio_async_out_i(30 downto 29);
    gt0_rxbufreset_i                             <= rx_data_vio_async_out_i(28);
    gt0_rxpmareset_i                             <= rx_data_vio_async_out_i(27);
    gt0_rxpolarity_i                             <= rx_data_vio_sync_out_i(31);
    gt0_ila_in_i(163 downto 162)                 <= gt0_rxchariscomma_i;
    gt0_ila_in_i(161 downto 160)                 <= gt0_rxcharisk_i;
    gt0_ila_in_i(159 downto 158)                 <= gt0_rxdisperr_i;
    gt0_ila_in_i(157 downto 156)                 <= gt0_rxnotintable_i;
    gt0_ila_in_i(155 downto 154)                 <= gt0_rxclkcorcnt_i;
    gt0_ila_in_i(153 downto 138)                 <= gt0_rxdata_i;
    gt0_ila_in_i(137 downto 135)                 <= gt0_rxbufstatus_i;
    gt0_ila_in_i(134 downto 127)                 <= gt0_error_count_i;
    gt0_ila_in_i(126)                            <= gt0_track_data_i;
    gt0_ila_in_i(125 downto 0)                   <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    gt0_channel_drp_vio_async_in_i(31)           <= gt0_drprdy_i;
    gt0_channel_drp_vio_async_in_i(30 downto 15) <= gt0_drpdo_i;
    gt0_channel_drp_vio_async_in_i(14 downto 0)  <= "000000000000000";
    gt0_channel_drp_vio_sync_in_i(31 downto 0)   <= "00000000000000000000000000000000";
    gt0_drpaddr_i                                <= channel_drp_vio_async_out_i(31 downto 23);
    gt0_drpdi_i                                  <= channel_drp_vio_async_out_i(22 downto 7);
    gt0_drpen_i                                  <= channel_drp_vio_async_out_i(6);
    gt0_drpwe_i                                  <= channel_drp_vio_async_out_i(5);
    gt0_common_drp_vio_async_in_i(31 downto 0)   <= "00000000000000000000000000000000";
    gt0_common_drp_vio_sync_in_i(31 downto 0)    <= "00000000000000000000000000000000";


    tx_data_vio_async_in_i              <=      gt0_tx_data_vio_async_in_i;

    tx_data_vio_sync_in_i               <=      gt0_tx_data_vio_sync_in_i;


    rx_data_vio_async_in_i              <=      gt0_rx_data_vio_async_in_i;

    rx_data_vio_sync_in_i               <=      gt0_rx_data_vio_sync_in_i;

    ila_in_i                            <=      gt0_ila_in_i;


    channel_drp_vio_async_in_i          <=      gt0_channel_drp_vio_async_in_i;

    channel_drp_vio_sync_in_i           <=      gt0_channel_drp_vio_sync_in_i;

    common_drp_vio_async_in_i <= (others => '0');
    common_drp_vio_sync_in_i  <= (others => '0');

end generate chipscope;

no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate

    -- assign resets for frame_gen modules
    gt0_tx_system_reset_c                        <= not gt0_txfsmresetdone_r2;

    -- assign resets for frame_check modules
    gt0_rx_system_reset_c                        <= not gt0_rxresetdone_r3;

    gttxreset_i                                  <= tied_to_ground_i;
    gtrxreset_i                                  <= tied_to_ground_i;
    user_tx_reset_i                              <= tied_to_ground_i;
    user_rx_reset_i                              <= tied_to_ground_i;
    gt0_loopback_i                               <= tied_to_ground_vec_i(2 downto 0);
    gt0_txpd_i                                   <= tied_to_ground_vec_i(1 downto 0);
    gt0_txchardispmode_i                         <= tied_to_ground_vec_i(1 downto 0);
    gt0_txchardispval_i                          <= tied_to_ground_vec_i(1 downto 0);
    gt0_txpolarity_i                             <= tied_to_ground_i;
    gt0_txelecidle_i                             <= tied_to_ground_i;
    gt0_rxpd_i                                   <= tied_to_ground_vec_i(1 downto 0);
    gt0_rxbufreset_i                             <= tied_to_ground_i;
    gt0_rxpmareset_i                             <= tied_to_ground_i;
    gt0_rxpolarity_i                             <= tied_to_ground_i;
    gt0_drpaddr_i                                <= tied_to_ground_vec_i(8 downto 0);
    gt0_drpdi_i                                  <= tied_to_ground_vec_i(15 downto 0);
    gt0_drpen_i                                  <= tied_to_ground_i;
    gt0_drpwe_i                                  <= tied_to_ground_i;


end generate no_chipscope;
end RTL;


